///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// Created by  : Prof. Quinn and Saumil Gogri
///////////////////////////////////////////////////////////////////////////

`include "base_test.sv"
`include "simple_random_test.sv"
`include "multiport_sequential_random_test.sv"
`include "short_packet_random_test.sv"
`include "medium_packet_random_test.sv"
`include "long_packet_random_test.sv"
`include "fixed_length_test.sv"
